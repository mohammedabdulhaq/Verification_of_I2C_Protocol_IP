class sequencer_0 extends uvm_sequencer#(sequence_item_0);
`uvm_object_utils(sequencer_0)

function new(string name = "sequencer_0", uvm_component parent = null);
        	super.new(name, parent);
        endfunction
function void build_phase(uvm_phase phase);
            super.build_phase(phase);
        endfunction

endclass